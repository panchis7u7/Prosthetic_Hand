module Seven_Segment_Display_Controller(
	input clk,
	input [11:0] data,
	output [3:0] select,
	output reg [7:0] lcd
);

always @(posedge clk)
begin
	
end

endmodule